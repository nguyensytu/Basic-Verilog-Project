module cpu (
    
);
    core core (clk, reset, inst, pc, data, data_valid);
    mem_map memory_map ();
endmodule