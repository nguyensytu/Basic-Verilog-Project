LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;
ENTITY tb_comparator IS
END tb_comparator;
ARCHITECTURE behavior OF tb_comparator IS 
    -- Component Declaration for the Unit Under Test (UUT)
    -- COMPONENT comparator
    -- PORT(
    --      clock : IN  std_logic;
    --      A : IN  std_logic_vector(7 downto 0);
    --      B : IN  std_logic_vector(7 downto 0);
    --      IAB : IN  std_logic;
    --      Output : OUT  std_logic
    --     );
    -- END COMPONENT;
   --Inputs
   signal clock : std_logic := '0';
   signal A : std_logic_vector(7 downto 0) := (others => '0');
   signal B : std_logic_vector(7 downto 0) := (others => '0');
   signal IAB : std_logic := '0';
 --Outputs
   signal Output : std_logic;
   -- Clock period definitions
   constant clock_period : time := 10 ns;
BEGIN
  -- Instantiate the Unit Under Test (UUT)
    uut: entity work.comparator 
    PORT MAP (
        clock => clock,
        A => A,
        B => B,
        IAB => IAB,
        Output => Output
    );
    -- Clock process definitions
    clock_process :process
    begin
        clock <= '0';
        wait for clock_period/2;
        clock <= '1';
        wait for clock_period/2;
    end process;
    -- Stimulus process
    stim_proc: process
    begin 
       -- hold reset state for 100 ns.
        wait for 100 ns; 
        A <= x"AA";
        B <= x"BB";
        wait for clock_period*10;
        B <= x"AA";
       -- insert stimulus here 
        wait;
    end process;
END;