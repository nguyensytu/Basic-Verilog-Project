module dma_priority (dma_if.PR dif, DmaControlIf.PR cif, DmaRegIf.PR rif);
    
endmodule