module uart_avalon #(
    parameter P = 0,
              EVEN_ODD = 0, // even  ~ 1, odd ~ 0
              W = 4,
              s = 1,
			  TIMER = 434
) (
    // Avalon interface
	input [1:0] address,
	input chipselect,
	input clk,
	input read,
	input reset_n,
	input write,
	input [31:0] writedata,
    output reg [31:0] readdata,
    // output
	input tdi,
    output wire tdo
);
// Signal declaration
    reg [31:0] data_tx, data_rx, status, control;
    reg [7+P:0] w_data; 
    wire [7+P:0] r_data;
    wire start, wr, rd, full_fifo_tx, empty_fifo_tx, full_fifo_rx, empty_fifo_rx, tx_tick, rx_tick;
    wire sum, parity;
// Submodule instance tx_fifo
    uart_tx_fifo #(.P(P), .W(W), .s(s), .TIMER(TIMER)) uart_tx_fifo (
        .clk(clk), .reset(~reset_n), .wr(wr), .start(start), .w_data(w_data), .full(full_fifo_tx), .empty(empty_fifo_tx), .tdo(tdo), .tx_tick(tx_tick)
    );
    single_cycle_tick start_cofigure (
        clk, ~reset_n, control[1], start
    );
    single_cycle_tick wr_configure (
        clk, ~reset_n, control[0], wr
    );
    assign sum = data_tx[0] + data_tx[1] + data_tx[2] + data_tx[3] + data_tx[4] + data_tx[5] + data_tx[6] + data_tx[7];
    assign parity = (EVEN_ODD) ? ~sum : sum;
    always @(*) begin
        if(P == 1)
            w_data = {parity, data_tx[7:0]};
        else    
            w_data = data_rx [7:0];
    end
// Submodule instance rx_fifo
    uart_rx_fifo #(.P(P), .W(W), .s(s), .TIMER(TIMER)) uart_rx_fifo (
        .clk(clk), .reset(~reset_n), .tdi(tdi), .rd(rd), .r_data(r_data), .empty(empty_fifo_rx), .full(full_fifo_rx), .rx_tick(rx_tick) 
    );
    single_cycle_tick rd_cofigure (
        clk, ~reset_n, control[2], rd
    );
// Avalon write/read
    always @(posedge clk or negedge reset_n) begin
        if(!reset_n) begin
            status [31:0] <= 32'b0;
            data_rx [31:0] <= 32'b0;
		end
        else begin
            status [31:6] <= 21'b0;
            data_rx [31:8+P] <= 21'b0; 
			status[5:0] <= {rx_tick, tx_tick, empty_fifo_rx, full_fifo_rx, empty_fifo_tx, full_fifo_tx};
            data_rx [7+P:0] <= r_data;
        end
    end
    always @ ( posedge clk or negedge reset_n )
	begin
		if ( reset_n == 1'b0 )
		begin
			data_tx <= 32'b0;
			control <= 32'b0;
			readdata <= 32'b0;
		end
		else if ( chipselect && write )
		begin
			case ( address )
				0 : data_tx <= writedata;
				3 : control <= writedata;
			endcase
		end
		else if ( chipselect && read )
		begin
			case ( address )
				0 : readdata <= data_tx;
                1 : readdata <= data_rx;
				2 : readdata <= status;
				3 : readdata <= control;
			endcase
		end
		else
		begin
			data_tx <= data_tx;
			control <= {control[31:3], rd, start, wr};
			readdata <= 32'b0;
		end
	end
endmodule